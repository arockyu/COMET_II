module RAM_256x16(
    input [7:0] addr,
    input [15:0] wdata,
    output [15:0] rdata,
    input ce,
    input clk,
    input we,
    input re);

    SB_RAM40_4K RAM_inst(
        .RDATA(rdata),
        .RADDR({3'b000,addr}),
        .RCLK(clk),
        .RCLKE(re&ce),
        .RE(re&ce),
        .WDATA(wdata),
        .WADDR({3'b000,addr}),
        .WCLK(clk),
        .WCLKE(we&ce),
        .WE(we&ce));
    defparam RAM_inst.READ_MODE =0;
    defparam RAM_inst.WRITE_MODE =0;

    defparam RAM_inst.INIT_1=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_2=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_3=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_4=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_5=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_6=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_7=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_8=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_9=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_A=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_B=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_C=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_D=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_E=
        256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam RAM_inst.INIT_F=
        256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule
