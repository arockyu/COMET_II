/************************************************************************
* Hex to 7-Seg decoder unit
*
*************************************************************************
* input [3:0] hex       : 1 digit hex(4-bit) input
* output [6:0] pat7seg : coded 7seg pattern output {g,f,e,d,c,b,a}
***************************************************************************
*  
* 
****************************************************************************/

module hexto7seg(
    input [3:0] hex,
    output [6:0] pat7seg);

    assign pat7seg = ( hex ==  4'h0 ) ? 7'b0111111 :
                     ( hex ==  4'h1 ) ? 7'b0000110 :     
                     ( hex ==  4'h2 ) ? 7'b1011011 :     
                     ( hex ==  4'h3 ) ? 7'b1001111 : 
                     ( hex ==  4'h4 ) ? 7'b1100110 : 
                     ( hex ==  4'h5 ) ? 7'b1101101 : 
                     ( hex ==  4'h6 ) ? 7'b1111101 : 
                     ( hex ==  4'h7 ) ? 7'b0000111 : 
                     ( hex ==  4'h8 ) ? 7'b1111111 : 
                     ( hex ==  4'h9 ) ? 7'b1101111 : 
                     ( hex ==  4'ha ) ? 7'b1110111 : 
                     ( hex ==  4'hb ) ? 7'b1111100 : 
                     ( hex ==  4'hc ) ? 7'b0111001 : 
                     ( hex ==  4'hd ) ? 7'b1011110 : 
                     ( hex ==  4'he ) ? 7'b1111001 : 
                     ( hex ==  4'hf ) ? 7'b1110001 : 7'b0000000; 
endmodule